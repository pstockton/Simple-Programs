`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// 64 x 64 Array Multiplier Test Bench
//
//  by: Patrick Stockton
//          
//
// 
//////////////////////////////////////////////////////////////////////////////////


module ArrayMult64x64_tb( );
    
    reg [63:0] A;
    reg [63:0] B;
    wire [127:0] Prod;
    
    ArrayMult64x64 UUT (.Prod(Prod), .A(A), .B(B));
    
    initial
    begin
        
        #100;
        
        // Reset A and B
        A = 16'h0000_0000_0000_0000; // A = 0
        B = 16'h0000_0000_0000_0000; // B = 0
        
        #20;
        // 2 * 8 = 16
        A = 16'h0000_0000_0000_0002; // A = 2
        B = 16'h0000_0000_0000_0008; // B = 8
        
        #20;
        // 10 * 32 = 320
        A = 16'h0000_0000_0000_000A; // A = 10
        B = 16'h0000_0000_0000_0020; // B = 32
        
        #20;
        // 256 * 512 = 131072
        A = 16'h0000_0000_0000_0100; // A = 256
        B = 16'h0000_0000_0000_0200; // B = 512
        
        #20;
        // 3000 * 55000
        A = 16'h0000_0000_0000_0BB8; // A = 3000
        B = 16'h0000_0000_0000_06D8; // B = 55000
      
    end
	
endmodule
