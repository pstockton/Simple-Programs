`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// 16-bit Carry Lookahead Adder Test Bench
//
// by: Patrick Stockton
//      
//
// 
//////////////////////////////////////////////////////////////////////////////////

module CLA16bit_tb( );
    reg [15:0] A, B;
    reg Cin;
    wire Cout, GG, PG;
    wire [15:0] S;
    
    CLA16bit UUT (.A(A), .B(B), .Cin(Cin), .S(S), .Cout(Cout), .GG(GG), .PG(PG));
        
    initial
    begin
        #100;
        A = 16'b0000000000000000;
        B = 16'b0000000000000000;
        Cin = 1'b0;
        
        #20;
        A = 8'b0000000000001111;
        B = 8'b0000000000000001;
        
        #20;
        B = 8'b0000000000000000;
        Cin = 1'b1;
        
        #20;
        Cin = 1'b0;
        A = 16'b1111111111111111;
        B = 16'b0000000000000001;
        
        #20;
        A = 16'b0101010101010101;
        B = 16'b1010101010101010;
        
        #20;
        Cin = 1'b1;       
    end
        
endmodule
