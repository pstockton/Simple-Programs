`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// 16-bit Ripple Carry Adder Test Bench
//
//	by: Patrick Stockton
// 
//////////////////////////////////////////////////////////////////////////////////


module RCA16bit_tb(  );

    reg [15:0] a, b;
    reg cin;
    wire [15:0] sum;
    wire cout;
    
    RCA16bit UUT (.sum(sum), .cout(cout), .a(a), .b(b), .cin(cin));
    
    initial
    begin
        a = 0;
        b = 0;
        cin = 0;
        
        #100;
        a = 16'b0000_0000_0000_1000;
        b = 16'b0000_0000_0000_0010;
        cin = 1'b0;
        
        #100;
        cin = 1'b1;
        
        #100;
        a = 16'b1000_0000_0000_0000;
        b = 16'b0000_0011_0000_0010;
        cin = 1'b0;
        
        #100;
        a = 16'b0000_0000_0100_1000;
        b = 16'b0000_0000_0000_1010;
        
        #100;
        a = 16'b0000_0000_0100_1000;
        b = 16'b1111_1111_1111_1111;
        
        #100;
        a = 16'b0000_0000_0000_0000;
        b = 16'b0000_0000_0000_0000;
                 
    end
	
endmodule
